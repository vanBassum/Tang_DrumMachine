module sine_rom(
    input  wire [7:0] addr,
    output reg  [9:0] data
);

    always @* begin
        case (addr)
            8'd0: data = 10'd512;
            8'd1: data = 10'd525;
            8'd2: data = 10'd537;
            8'd3: data = 10'd550;
            8'd4: data = 10'd562;
            8'd5: data = 10'd575;
            8'd6: data = 10'd587;
            8'd7: data = 10'd599;
            8'd8: data = 10'd612;
            8'd9: data = 10'd624;
            8'd10: data = 10'd636;
            8'd11: data = 10'd648;
            8'd12: data = 10'd660;
            8'd13: data = 10'd672;
            8'd14: data = 10'd684;
            8'd15: data = 10'd696;
            8'd16: data = 10'd708;
            8'd17: data = 10'd719;
            8'd18: data = 10'd730;
            8'd19: data = 10'd742;
            8'd20: data = 10'd753;
            8'd21: data = 10'd764;
            8'd22: data = 10'd775;
            8'd23: data = 10'd785;
            8'd24: data = 10'd796;
            8'd25: data = 10'd806;
            8'd26: data = 10'd816;
            8'd27: data = 10'd826;
            8'd28: data = 10'd836;
            8'd29: data = 10'd846;
            8'd30: data = 10'd855;
            8'd31: data = 10'd864;
            8'd32: data = 10'd873;
            8'd33: data = 10'd882;
            8'd34: data = 10'd891;
            8'd35: data = 10'd899;
            8'd36: data = 10'd907;
            8'd37: data = 10'd915;
            8'd38: data = 10'd922;
            8'd39: data = 10'd930;
            8'd40: data = 10'd937;
            8'd41: data = 10'd944;
            8'd42: data = 10'd950;
            8'd43: data = 10'd957;
            8'd44: data = 10'd963;
            8'd45: data = 10'd968;
            8'd46: data = 10'd974;
            8'd47: data = 10'd979;
            8'd48: data = 10'd984;
            8'd49: data = 10'd989;
            8'd50: data = 10'd993;
            8'd51: data = 10'd997;
            8'd52: data = 10'd1001;
            8'd53: data = 10'd1004;
            8'd54: data = 10'd1008;
            8'd55: data = 10'd1011;
            8'd56: data = 10'd1013;
            8'd57: data = 10'd1015;
            8'd58: data = 10'd1017;
            8'd59: data = 10'd1019;
            8'd60: data = 10'd1021;
            8'd61: data = 10'd1022;
            8'd62: data = 10'd1022;
            8'd63: data = 10'd1023;
            8'd64: data = 10'd1023;
            8'd65: data = 10'd1023;
            8'd66: data = 10'd1022;
            8'd67: data = 10'd1022;
            8'd68: data = 10'd1021;
            8'd69: data = 10'd1019;
            8'd70: data = 10'd1017;
            8'd71: data = 10'd1015;
            8'd72: data = 10'd1013;
            8'd73: data = 10'd1011;
            8'd74: data = 10'd1008;
            8'd75: data = 10'd1004;
            8'd76: data = 10'd1001;
            8'd77: data = 10'd997;
            8'd78: data = 10'd993;
            8'd79: data = 10'd989;
            8'd80: data = 10'd984;
            8'd81: data = 10'd979;
            8'd82: data = 10'd974;
            8'd83: data = 10'd968;
            8'd84: data = 10'd963;
            8'd85: data = 10'd957;
            8'd86: data = 10'd950;
            8'd87: data = 10'd944;
            8'd88: data = 10'd937;
            8'd89: data = 10'd930;
            8'd90: data = 10'd922;
            8'd91: data = 10'd915;
            8'd92: data = 10'd907;
            8'd93: data = 10'd899;
            8'd94: data = 10'd891;
            8'd95: data = 10'd882;
            8'd96: data = 10'd873;
            8'd97: data = 10'd864;
            8'd98: data = 10'd855;
            8'd99: data = 10'd846;
            8'd100: data = 10'd836;
            8'd101: data = 10'd826;
            8'd102: data = 10'd816;
            8'd103: data = 10'd806;
            8'd104: data = 10'd796;
            8'd105: data = 10'd785;
            8'd106: data = 10'd775;
            8'd107: data = 10'd764;
            8'd108: data = 10'd753;
            8'd109: data = 10'd742;
            8'd110: data = 10'd730;
            8'd111: data = 10'd719;
            8'd112: data = 10'd708;
            8'd113: data = 10'd696;
            8'd114: data = 10'd684;
            8'd115: data = 10'd672;
            8'd116: data = 10'd660;
            8'd117: data = 10'd648;
            8'd118: data = 10'd636;
            8'd119: data = 10'd624;
            8'd120: data = 10'd612;
            8'd121: data = 10'd599;
            8'd122: data = 10'd587;
            8'd123: data = 10'd575;
            8'd124: data = 10'd562;
            8'd125: data = 10'd550;
            8'd126: data = 10'd537;
            8'd127: data = 10'd525;
            8'd128: data = 10'd512;
            8'd129: data = 10'd499;
            8'd130: data = 10'd487;
            8'd131: data = 10'd474;
            8'd132: data = 10'd462;
            8'd133: data = 10'd449;
            8'd134: data = 10'd437;
            8'd135: data = 10'd425;
            8'd136: data = 10'd412;
            8'd137: data = 10'd400;
            8'd138: data = 10'd388;
            8'd139: data = 10'd376;
            8'd140: data = 10'd364;
            8'd141: data = 10'd352;
            8'd142: data = 10'd340;
            8'd143: data = 10'd328;
            8'd144: data = 10'd316;
            8'd145: data = 10'd305;
            8'd146: data = 10'd294;
            8'd147: data = 10'd282;
            8'd148: data = 10'd271;
            8'd149: data = 10'd260;
            8'd150: data = 10'd249;
            8'd151: data = 10'd239;
            8'd152: data = 10'd228;
            8'd153: data = 10'd218;
            8'd154: data = 10'd208;
            8'd155: data = 10'd198;
            8'd156: data = 10'd188;
            8'd157: data = 10'd178;
            8'd158: data = 10'd169;
            8'd159: data = 10'd160;
            8'd160: data = 10'd151;
            8'd161: data = 10'd142;
            8'd162: data = 10'd133;
            8'd163: data = 10'd125;
            8'd164: data = 10'd117;
            8'd165: data = 10'd109;
            8'd166: data = 10'd102;
            8'd167: data = 10'd94;
            8'd168: data = 10'd87;
            8'd169: data = 10'd80;
            8'd170: data = 10'd74;
            8'd171: data = 10'd67;
            8'd172: data = 10'd61;
            8'd173: data = 10'd56;
            8'd174: data = 10'd50;
            8'd175: data = 10'd45;
            8'd176: data = 10'd40;
            8'd177: data = 10'd35;
            8'd178: data = 10'd31;
            8'd179: data = 10'd27;
            8'd180: data = 10'd23;
            8'd181: data = 10'd20;
            8'd182: data = 10'd16;
            8'd183: data = 10'd13;
            8'd184: data = 10'd11;
            8'd185: data = 10'd9;
            8'd186: data = 10'd7;
            8'd187: data = 10'd5;
            8'd188: data = 10'd3;
            8'd189: data = 10'd2;
            8'd190: data = 10'd2;
            8'd191: data = 10'd1;
            8'd192: data = 10'd1;
            8'd193: data = 10'd1;
            8'd194: data = 10'd2;
            8'd195: data = 10'd2;
            8'd196: data = 10'd3;
            8'd197: data = 10'd5;
            8'd198: data = 10'd7;
            8'd199: data = 10'd9;
            8'd200: data = 10'd11;
            8'd201: data = 10'd13;
            8'd202: data = 10'd16;
            8'd203: data = 10'd20;
            8'd204: data = 10'd23;
            8'd205: data = 10'd27;
            8'd206: data = 10'd31;
            8'd207: data = 10'd35;
            8'd208: data = 10'd40;
            8'd209: data = 10'd45;
            8'd210: data = 10'd50;
            8'd211: data = 10'd56;
            8'd212: data = 10'd61;
            8'd213: data = 10'd67;
            8'd214: data = 10'd74;
            8'd215: data = 10'd80;
            8'd216: data = 10'd87;
            8'd217: data = 10'd94;
            8'd218: data = 10'd102;
            8'd219: data = 10'd109;
            8'd220: data = 10'd117;
            8'd221: data = 10'd125;
            8'd222: data = 10'd133;
            8'd223: data = 10'd142;
            8'd224: data = 10'd151;
            8'd225: data = 10'd160;
            8'd226: data = 10'd169;
            8'd227: data = 10'd178;
            8'd228: data = 10'd188;
            8'd229: data = 10'd198;
            8'd230: data = 10'd208;
            8'd231: data = 10'd218;
            8'd232: data = 10'd228;
            8'd233: data = 10'd239;
            8'd234: data = 10'd249;
            8'd235: data = 10'd260;
            8'd236: data = 10'd271;
            8'd237: data = 10'd282;
            8'd238: data = 10'd294;
            8'd239: data = 10'd305;
            8'd240: data = 10'd316;
            8'd241: data = 10'd328;
            8'd242: data = 10'd340;
            8'd243: data = 10'd352;
            8'd244: data = 10'd364;
            8'd245: data = 10'd376;
            8'd246: data = 10'd388;
            8'd247: data = 10'd400;
            8'd248: data = 10'd412;
            8'd249: data = 10'd425;
            8'd250: data = 10'd437;
            8'd251: data = 10'd449;
            8'd252: data = 10'd462;
            8'd253: data = 10'd474;
            8'd254: data = 10'd487;
            8'd255: data = 10'd499;
            default: data = 10'd512;
        endcase
    end

endmodule
